/*************************************************************************
 > File Name: test.v
 > Author: Darphee
  Last Modified: 2023年06月17日 星期六 00时16分18秒
 ************************************************************************/


module



endmodule

